library verilog;
use verilog.vl_types.all;
entity Master_vlg_vec_tst is
end Master_vlg_vec_tst;
